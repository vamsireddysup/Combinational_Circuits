module Nto1_mux(#parameter N=2)(
	input bit [N-1:0][3:0]ip,
	input bit [$clog2(N)-1:0]sel,
	output bit [3:0]out
	);
	x



endmodule:Nto1_mux
