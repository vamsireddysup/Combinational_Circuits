module check

//check to commit
endmodule:check
