module check


endmodule:check
